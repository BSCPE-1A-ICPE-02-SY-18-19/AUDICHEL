CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 12 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 101 143 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
43530.4 0
0
2 +V
167 251 75 0 1 3
0 17
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7876 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 876 53 0 18 19
10 9 8 7 6 5 4 3 18 19
0 1 0 0 0 1 1 2 2
0
0 0 21088 0
8 YELLOWCC
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
6369 0 0
2
43530.3 0
0
9 2-In AND~
219 524 68 0 3 22
0 15 14 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9172 0 0
2
43530.3 0
0
9 2-In AND~
219 406 71 0 3 22
0 10 11 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7100 0 0
2
43530.3 0
0
6 74LS48
188 736 126 0 14 29
0 12 14 11 10 20 21 3 4 5
6 7 8 9 22
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
3820 0 0
2
43530.3 0
0
6 74112~
219 576 215 0 7 32
0 17 13 16 13 17 23 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
7678 0 0
2
43530.3 0
0
6 74112~
219 456 219 0 7 32
0 17 15 16 15 17 24 14
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
961 0 0
2
43530.3 0
0
6 74112~
219 342 220 0 7 32
0 17 10 16 10 17 25 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3178 0 0
2
43530.3 0
0
6 74112~
219 227 222 0 7 32
0 17 2 16 2 17 26 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3409 0 0
2
43530.3 0
0
7 Pulser~
4 99 275 0 10 12
0 27 28 29 16 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3951 0 0
2
43530.3 0
0
37
1 0 2 0 0 4224 0 1 0 0 2 3
113 143
187 143
187 186
4 2 2 0 0 0 0 10 10 0 0 4
203 204
187 204
187 186
203 186
7 7 3 0 0 8320 0 6 3 0 0 3
768 90
768 89
891 89
8 6 4 0 0 4224 0 6 3 0 0 3
768 99
885 99
885 89
9 5 5 0 0 4224 0 6 3 0 0 3
768 108
879 108
879 89
10 4 6 0 0 4224 0 6 3 0 0 3
768 117
873 117
873 89
11 3 7 0 0 4224 0 6 3 0 0 3
768 126
867 126
867 89
12 2 8 0 0 4224 0 6 3 0 0 3
768 135
861 135
861 89
13 1 9 0 0 4224 0 6 3 0 0 3
768 144
855 144
855 89
4 0 10 0 0 4224 0 6 0 0 25 3
704 117
275 117
275 184
3 0 11 0 0 4224 0 6 0 0 18 2
704 108
366 108
1 7 12 0 0 4224 0 6 7 0 0 3
704 90
600 90
600 179
2 0 13 0 0 4096 0 7 0 0 14 2
552 179
545 179
4 3 13 0 0 8320 0 7 4 0 0 3
552 197
545 197
545 68
2 0 14 0 0 4224 0 6 0 0 17 2
704 99
480 99
1 3 15 0 0 4096 0 4 5 0 0 3
500 59
427 59
427 71
7 2 14 0 0 0 0 8 4 0 0 3
480 183
480 77
500 77
7 2 11 0 0 0 0 9 5 0 0 3
366 184
366 80
382 80
2 0 15 0 0 0 0 8 0 0 20 3
432 183
432 151
427 151
3 4 15 0 0 4224 0 5 8 0 0 5
427 71
427 151
412 151
412 201
432 201
3 0 16 0 0 4096 0 8 0 0 37 2
426 192
426 275
3 0 16 0 0 0 0 9 0 0 37 2
312 193
312 275
0 1 10 0 0 0 0 0 5 24 0 3
299 185
299 62
382 62
4 0 10 0 0 0 0 9 0 0 25 3
318 202
299 202
299 184
7 2 10 0 0 0 0 10 9 0 0 3
251 186
251 184
318 184
1 0 17 0 0 4096 0 2 0 0 32 2
251 84
251 123
0 0 17 0 0 4096 0 0 0 32 35 2
287 123
287 242
0 0 17 0 0 0 0 0 0 32 35 2
399 123
399 242
0 0 17 0 0 0 0 0 0 32 35 2
497 123
497 242
1 0 17 0 0 0 0 8 0 0 32 2
456 156
456 123
1 0 17 0 0 0 0 9 0 0 32 2
342 157
342 123
1 1 17 0 0 8320 0 10 7 0 0 4
227 159
227 123
576 123
576 152
5 0 17 0 0 0 0 8 0 0 35 2
456 231
456 242
5 0 17 0 0 0 0 9 0 0 35 2
342 232
342 242
5 5 17 0 0 16 0 10 7 0 0 4
227 234
227 242
576 242
576 227
3 0 16 0 0 0 0 10 0 0 37 2
197 195
197 275
4 3 16 0 0 4224 0 11 7 0 0 4
129 275
510 275
510 188
546 188
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
